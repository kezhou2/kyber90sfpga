module mem_gen5 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 12;
input clk;
input [5:0] addr;
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= 12'd2285;
1: data <= 12'd1701;
2: data <= 12'd1275;
3: data <= 12'd75;
4: data <= 12'd1571;
5: data <= 12'd1659;
6: data <= 12'd1860;
7: data <= 12'd1676;
8: data <= 12'd1861;
9: data <= 12'd2851;
10: data <= 12'd951;
11: data <= 12'd2210;
12: data <= 12'd130;
13: data <= 12'd2945;
14: data <= 12'd1544;
15: data <= 12'd3224;
16: data <= 12'd3127;
17: data <= 12'd2338;
18: data <= 12'd725;
19: data <= 12'd2980;
20: data <= 12'd2721;
21: data <= 12'd1335;
22: data <= 12'd666;
23: data <= 12'd235;
24: data <= 12'd3147;
25: data <= 12'd2535;
26: data <= 12'd2499;
27: data <= 12'd147;
28: data <= 12'd2946;
29: data <= 12'd2719;
30: data <= 12'd2314;
31: data <= 12'd2486;
32: data <= 12'd1517;
33: data <= 12'd1460;
34: data <= 12'd1065;
35: data <= 12'd3000;
36: data <= 12'd2918;
37: data <= 12'd3109;
38: data <= 12'd1162;
39: data <= 12'd460;
40: data <= 12'd1202;
41: data <= 12'd854;
42: data <= 12'd1421;
43: data <= 12'd1846;
44: data <= 12'd1871;
45: data <= 12'd1285;
46: data <= 12'd1838;
47: data <= 12'd2458;
48: data <= 12'd1907;
49: data <= 12'd308;
50: data <= 12'd2368;
51: data <= 12'd2685;
52: data <= 12'd2312;
53: data <= 12'd136;
54: data <= 12'd8;
55: data <= 12'd2742;
56: data <= 12'd2707;
57: data <= 12'd1530;
58: data <= 12'd90;
59: data <= 12'd2551;
60: data <= 12'd1325;
61: data <= 12'd2232;
62: data <= 12'd2677;
63: data <= 12'd2899;
    default : data <= 0;
    endcase
end
endmodule
