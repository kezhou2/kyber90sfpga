module mem_gen1 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 12;
input clk;
input [5:0] addr;
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= 12'd2285;
1: data <= 12'd2226;
2: data <= 12'd1223;
3: data <= 12'd817;
4: data <= 12'd573;
5: data <= 12'd3083;
6: data <= 12'd2476;
7: data <= 12'd2144;
8: data <= 12'd3158;
9: data <= 12'd422;
10: data <= 12'd516;
11: data <= 12'd2114;
12: data <= 12'd2648;
13: data <= 12'd1739;
14: data <= 12'd2931;
15: data <= 12'd3221;
16: data <= 12'd1493;
17: data <= 12'd2078;
18: data <= 12'd2036;
19: data <= 12'd1322;
20: data <= 12'd2500;
21: data <= 12'd2552;
22: data <= 12'd107;
23: data <= 12'd1819;
24: data <= 12'd962;
25: data <= 12'd3038;
26: data <= 12'd1711;
27: data <= 12'd2455;
28: data <= 12'd1787;
29: data <= 12'd418;
30: data <= 12'd448;
31: data <= 12'd958;
32: data <= 12'd2970;
33: data <= 12'd555;
34: data <= 12'd2777;
35: data <= 12'd603;
36: data <= 12'd264;
37: data <= 12'd1159;
38: data <= 12'd3058;
39: data <= 12'd2051;
40: data <= 12'd1577;
41: data <= 12'd177;
42: data <= 12'd3009;
43: data <= 12'd1218;
44: data <= 12'd732;
45: data <= 12'd2457;
46: data <= 12'd1821;
47: data <= 12'd996;
48: data <= 12'd287;
49: data <= 12'd1550;
50: data <= 12'd3047;
51: data <= 12'd1864;
52: data <= 12'd1727;
53: data <= 12'd2727;
54: data <= 12'd3082;
55: data <= 12'd2459;
56: data <= 12'd1855;
57: data <= 12'd1574;
58: data <= 12'd126;
59: data <= 12'd2142;
60: data <= 12'd3124;
61: data <= 12'd3173;
62: data <= 12'd677;
63: data <= 12'd1522;
    default : data <= 0;
    endcase
end
endmodule
