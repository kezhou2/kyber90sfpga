////////////////////////////////////////////////////////////////////////////////
//
// Hung Technologies
//
// Filename     : mux_xx1.v
// Description  : .
//
// Author       : hungnt@HW-NTHUNG
// Created On   : Thu Nov 08 10:51:52 2018
// History (Date, Changed By)
//
////////////////////////////////////////////////////////////////////////////////

module mux_xx2
    (
     a,
     b,
     c,
     d,
     s,
     o
     );

////////////////////////////////////////////////////////////////////////////////
// Parameter declarations

parameter WIDTH = 1;

////////////////////////////////////////////////////////////////////////////////
// Port declarations

////////////////////////////////////////////////////////////////////////////////
// Output declarations

input     s;
input [WIDTH-1:0] a,b,c,d;

output [WIDTH-1:0] o;

////////////////////////////////////////////////////////////////////////////////
// Local logic and instantiation

always @(*) case(sel)
	2'h 0 : o = a;
	2'h 1 : o = b;
	2'h 2 : o = c;
	default : o = d;
endcase

endmodule 
