module mem_gen5 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 12;
input clk;
input [6:0] addr;
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= 12'd2285;
1: data <= 12'd2044;
2: data <= 12'd271;
3: data <= 12'd1676;
4: data <= 12'd1017;
5: data <= 12'd2371;
6: data <= 12'd1544;
7: data <= 12'd778;
8: data <= 12'd2367;
9: data <= 12'd1335;
10: data <= 12'd677;
11: data <= 12'd1251;
12: data <= 12'd2946;
13: data <= 12'd2459;
14: data <= 12'd2813;
15: data <= 12'd3000;
16: data <= 12'd287;
17: data <= 12'd2512;
18: data <= 12'd1421;
19: data <= 12'd177;
20: data <= 12'd1758;
21: data <= 12'd308;
22: data <= 12'd2777;
23: data <= 12'd1119;
24: data <= 12'd2707;
25: data <= 12'd2455;
26: data <= 12'd2604;
27: data <= 12'd2899;
28: data <= 12'd2500;
29: data <= 12'd794;
30: data <= 12'd3203;
31: data <= 12'd1739;
32: data <= 12'd1812;
33: data <= 12'd1465;
34: data <= 12'd2476;
35: data <= 12'd2869;
36: data <= 12'd2597;
37: data <= 12'd1701;
38: data <= 12'd1491;
39: data <= 12'd2170;
40: data <= 12'd1861;
41: data <= 12'd3193;
42: data <= 12'd2881;
43: data <= 12'd3224;
44: data <= 12'd2004;
45: data <= 12'd1510;
46: data <= 12'd666;
47: data <= 12'd3173;
48: data <= 12'd1836;
49: data <= 12'd2719;
50: data <= 12'd3082;
51: data <= 12'd2907;
52: data <= 12'd2918;
53: data <= 12'd996;
54: data <= 12'd2106;
55: data <= 12'd1846;
56: data <= 12'd1577;
57: data <= 12'd1670;
58: data <= 12'd2368;
59: data <= 12'd555;
60: data <= 12'd3199;
61: data <= 12'd1530;
62: data <= 12'd1711;
63: data <= 12'd349;
64: data <= 12'd758;
65: data <= 12'd1322;
66: data <= 12'd830;
67: data <= 12'd1755;
68: data <= 12'd2648;
69: data <= 12'd1869;
70: data <= 12'd282;
71: data <= 12'd3083;
72: data <= 12'd2127;
73: data <= 12'd2111;
74: data <= 12'd1275;
75: data <= 12'd871;
76: data <= 12'd3065;
77: data <= 12'd2851;
78: data <= 12'd3321;
79: data <= 12'd2911;
80: data <= 12'd3127;
81: data <= 12'd1097;
82: data <= 12'd3222;
83: data <= 12'd235;
84: data <= 12'd3124;
85: data <= 12'd108;
86: data <= 12'd2314;
87: data <= 12'd2727;
88: data <= 12'd171;
89: data <= 12'd3109;
90: data <= 12'd1821;
91: data <= 12'd1103;
92: data <= 12'd1871;
93: data <= 12'd2051;
94: data <= 12'd1469;
95: data <= 12'd2685;
96: data <= 12'd2970;
97: data <= 12'd384;
98: data <= 12'd90;
99: data <= 12'd3038;
100: data <= 12'd608;
101: data <= 12'd1807;
102: data <= 12'd2036;
103: data <= 12'd3182;
104: data <= 12'd1474;
105: data <= 12'd2114;
106: data <= 12'd2264;
107: data <= 12'd1779;
108: data <= 12'd573;
109: data <= 12'd2475;
110: data <= 12'd320;
111: data <= 12'd75;
112: data <= 12'd1422;
113: data <= 12'd2726;
114: data <= 12'd951;
115: data <= 12'd587;
116: data <= 12'd1542;
117: data <= 12'd2338;
118: data <= 12'd652;
119: data <= 12'd777;
120: data <= 12'd3147;
121: data <= 12'd2142;
122: data <= 12'd398;
123: data <= 12'd2486;
124: data <= 12'd1727;
125: data <= 12'd1185;
126: data <= 12'd1162;
127: data <= 12'd2457;
    default : data <= 0;
    endcase
end
endmodule
