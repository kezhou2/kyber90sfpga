module polyunit(
    clk,
    rst,
    
)