module mem_gen6 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 7*4;
input clk;
input [6:0] addr;//127
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= {7'd1,7'd9,7'd0,7'd0};
1: data <= {7'd3,7'd11,7'd0,7'd0};
2: data <= {7'd5,7'd13,7'd0,7'd0};
3: data <= {7'd7,7'd15,7'd0,7'd0};
4: data <= {7'd17,7'd25,7'd0,7'd0};
5: data <= {7'd19,7'd27,7'd0,7'd0};
6: data <= {7'd21,7'd29,7'd0,7'd0};
7: data <= {7'd23,7'd31,7'd0,7'd0};
8: data <= {7'd33,7'd41,7'd0,7'd0};
9: data <= {7'd35,7'd43,7'd0,7'd0};
10: data <= {7'd37,7'd45,7'd0,7'd0};
11: data <= {7'd39,7'd47,7'd0,7'd0};
12: data <= {7'd49,7'd57,7'd0,7'd0};
13: data <= {7'd51,7'd59,7'd0,7'd0};
14: data <= {7'd53,7'd61,7'd0,7'd0};
15: data <= {7'd55,7'd63,7'd0,7'd0};
16: data <= {7'd65,7'd73,7'd0,7'd0};
17: data <= {7'd67,7'd75,7'd0,7'd0};
18: data <= {7'd69,7'd77,7'd0,7'd0};
19: data <= {7'd71,7'd79,7'd0,7'd0};
20: data <= {7'd81,7'd89,7'd0,7'd0};
21: data <= {7'd83,7'd91,7'd0,7'd0};
22: data <= {7'd85,7'd93,7'd0,7'd0};
23: data <= {7'd87,7'd95,7'd0,7'd0};
24: data <= {7'd97,7'd105,7'd0,7'd0};
25: data <= {7'd99,7'd107,7'd0,7'd0};
26: data <= {7'd101,7'd109,7'd0,7'd0};
27: data <= {7'd103,7'd111,7'd0,7'd0};
28: data <= {7'd113,7'd121,7'd0,7'd0};
29: data <= {7'd115,7'd123,7'd0,7'd0};
30: data <= {7'd117,7'd125,7'd0,7'd0};
31: data <= {7'd119,7'd127,7'd0,7'd0};
32: data <= {7'd4,7'd4,7'd66,7'd2};
33: data <= {7'd68,7'd68,7'd98,7'd34};
34: data <= {7'd36,7'd36,7'd82,7'd18};
35: data <= {7'd100,7'd100,7'd114,7'd50};
36: data <= {7'd4,7'd4,7'd66,7'd2};
37: data <= {7'd68,7'd68,7'd98,7'd34};
38: data <= {7'd36,7'd36,7'd82,7'd18};
39: data <= {7'd100,7'd100,7'd114,7'd50};
40: data <= {7'd20,7'd20,7'd74,7'd10};
41: data <= {7'd84,7'd84,7'd106,7'd42};
42: data <= {7'd52,7'd52,7'd90,7'd26};
43: data <= {7'd116,7'd116,7'd122,7'd58};
44: data <= {7'd20,7'd20,7'd74,7'd10};
45: data <= {7'd84,7'd84,7'd106,7'd42};
46: data <= {7'd52,7'd52,7'd90,7'd26};
47: data <= {7'd116,7'd116,7'd122,7'd58};
48: data <= {7'd12,7'd12,7'd70,7'd6};
49: data <= {7'd76,7'd76,7'd102,7'd38};
50: data <= {7'd44,7'd44,7'd86,7'd22};
51: data <= {7'd108,7'd108,7'd118,7'd54};
52: data <= {7'd12,7'd12,7'd70,7'd6};
53: data <= {7'd76,7'd76,7'd102,7'd38};
54: data <= {7'd44,7'd44,7'd86,7'd22};
55: data <= {7'd108,7'd108,7'd118,7'd54};
56: data <= {7'd28,7'd28,7'd78,7'd14};
57: data <= {7'd92,7'd92,7'd110,7'd46};
58: data <= {7'd60,7'd60,7'd94,7'd30};
59: data <= {7'd124,7'd124,7'd126,7'd62};
60: data <= {7'd28,7'd28,7'd78,7'd14};
61: data <= {7'd92,7'd92,7'd110,7'd46};
62: data <= {7'd60,7'd60,7'd94,7'd30};
63: data <= {7'd124,7'd124,7'd126,7'd62};
64: data <= {7'd16,7'd16,7'd72,7'd8};
65: data <= {7'd80,7'd80,7'd104,7'd40};
66: data <= {7'd48,7'd48,7'd88,7'd24};
67: data <= {7'd112,7'd112,7'd120,7'd56};
68: data <= {7'd16,7'd16,7'd72,7'd8};
69: data <= {7'd80,7'd80,7'd104,7'd40};
70: data <= {7'd48,7'd48,7'd88,7'd24};
71: data <= {7'd112,7'd112,7'd120,7'd56};
72: data <= {7'd16,7'd16,7'd72,7'd8};
73: data <= {7'd80,7'd80,7'd104,7'd40};
74: data <= {7'd48,7'd48,7'd88,7'd24};
75: data <= {7'd112,7'd112,7'd120,7'd56};
76: data <= {7'd16,7'd16,7'd72,7'd8};
77: data <= {7'd80,7'd80,7'd104,7'd40};
78: data <= {7'd48,7'd48,7'd88,7'd24};
79: data <= {7'd112,7'd112,7'd120,7'd56};
80: data <= {7'd16,7'd16,7'd72,7'd8};
81: data <= {7'd80,7'd80,7'd104,7'd40};
82: data <= {7'd48,7'd48,7'd88,7'd24};
83: data <= {7'd112,7'd112,7'd120,7'd56};
84: data <= {7'd16,7'd16,7'd72,7'd8};
85: data <= {7'd80,7'd80,7'd104,7'd40};
86: data <= {7'd48,7'd48,7'd88,7'd24};
87: data <= {7'd112,7'd112,7'd120,7'd56};
88: data <= {7'd16,7'd16,7'd72,7'd8};
89: data <= {7'd80,7'd80,7'd104,7'd40};
90: data <= {7'd48,7'd48,7'd88,7'd24};
91: data <= {7'd112,7'd112,7'd120,7'd56};
92: data <= {7'd16,7'd16,7'd72,7'd8};
93: data <= {7'd80,7'd80,7'd104,7'd40};
94: data <= {7'd48,7'd48,7'd88,7'd24};
95: data <= {7'd112,7'd112,7'd120,7'd56};
96: data <= {7'd64,7'd64,7'd96,7'd32};
97: data <= {7'd64,7'd64,7'd96,7'd32};
98: data <= {7'd64,7'd64,7'd96,7'd32};
99: data <= {7'd64,7'd64,7'd96,7'd32};
100: data <= {7'd64,7'd64,7'd96,7'd32};
101: data <= {7'd64,7'd64,7'd96,7'd32};
102: data <= {7'd64,7'd64,7'd96,7'd32};
103: data <= {7'd64,7'd64,7'd96,7'd32};
104: data <= {7'd64,7'd64,7'd96,7'd32};
105: data <= {7'd64,7'd64,7'd96,7'd32};
106: data <= {7'd64,7'd64,7'd96,7'd32};
107: data <= {7'd64,7'd64,7'd96,7'd32};
108: data <= {7'd64,7'd64,7'd96,7'd32};
109: data <= {7'd64,7'd64,7'd96,7'd32};
110: data <= {7'd64,7'd64,7'd96,7'd32};
111: data <= {7'd64,7'd64,7'd96,7'd32};
112: data <= {7'd64,7'd64,7'd96,7'd32};
113: data <= {7'd64,7'd64,7'd96,7'd32};
114: data <= {7'd64,7'd64,7'd96,7'd32};
115: data <= {7'd64,7'd64,7'd96,7'd32};
116: data <= {7'd64,7'd64,7'd96,7'd32};
117: data <= {7'd64,7'd64,7'd96,7'd32};
118: data <= {7'd64,7'd64,7'd96,7'd32};
119: data <= {7'd64,7'd64,7'd96,7'd32};
120: data <= {7'd64,7'd64,7'd96,7'd32};
121: data <= {7'd64,7'd64,7'd96,7'd32};
122: data <= {7'd64,7'd64,7'd96,7'd32};
123: data <= {7'd64,7'd64,7'd96,7'd32};
124: data <= {7'd64,7'd64,7'd96,7'd32};
125: data <= {7'd64,7'd64,7'd96,7'd32};
126: data <= {7'd64,7'd64,7'd96,7'd32};
127: data <= {7'd64,7'd64,7'd96,7'd32};
    default : data <= 0;
    endcase
end
endmodule
