module mem_gen3 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 5;
input clk;
input [6:0] addr;
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= 5'd0;
1: data <= 5'd8;
2: data <= 5'd16;
3: data <= 5'd24;
4: data <= 5'd1;
5: data <= 5'd9;
6: data <= 5'd17;
7: data <= 5'd25;
8: data <= 5'd2;
9: data <= 5'd10;
10: data <= 5'd18;
11: data <= 5'd26;
12: data <= 5'd3;
13: data <= 5'd11;
14: data <= 5'd19;
15: data <= 5'd27;
16: data <= 5'd4;
17: data <= 5'd12;
18: data <= 5'd20;
19: data <= 5'd28;
20: data <= 5'd5;
21: data <= 5'd13;
22: data <= 5'd21;
23: data <= 5'd29;
24: data <= 5'd6;
25: data <= 5'd14;
26: data <= 5'd22;
27: data <= 5'd30;
28: data <= 5'd7;
29: data <= 5'd15;
30: data <= 5'd23;
31: data <= 5'd31;
32: data <= 5'd0;
33: data <= 5'd2;
34: data <= 5'd4;
35: data <= 5'd6;
36: data <= 5'd1;
37: data <= 5'd3;
38: data <= 5'd5;
39: data <= 5'd7;
40: data <= 5'd8;
41: data <= 5'd10;
42: data <= 5'd12;
43: data <= 5'd14;
44: data <= 5'd9;
45: data <= 5'd11;
46: data <= 5'd13;
47: data <= 5'd15;
48: data <= 5'd16;
49: data <= 5'd18;
50: data <= 5'd20;
51: data <= 5'd22;
52: data <= 5'd17;
53: data <= 5'd19;
54: data <= 5'd21;
55: data <= 5'd23;
56: data <= 5'd24;
57: data <= 5'd26;
58: data <= 5'd28;
59: data <= 5'd30;
60: data <= 5'd25;
61: data <= 5'd27;
62: data <= 5'd29;
63: data <= 5'd31;
64: data <= 5'd0;
65: data <= 5'd1;
66: data <= 5'd2;
67: data <= 5'd3;
68: data <= 5'd4;
69: data <= 5'd5;
70: data <= 5'd6;
71: data <= 5'd7;
72: data <= 5'd8;
73: data <= 5'd9;
74: data <= 5'd10;
75: data <= 5'd11;
76: data <= 5'd12;
77: data <= 5'd13;
78: data <= 5'd14;
79: data <= 5'd15;
80: data <= 5'd16;
81: data <= 5'd17;
82: data <= 5'd18;
83: data <= 5'd19;
84: data <= 5'd20;
85: data <= 5'd21;
86: data <= 5'd22;
87: data <= 5'd23;
88: data <= 5'd24;
89: data <= 5'd25;
90: data <= 5'd26;
91: data <= 5'd27;
92: data <= 5'd28;
93: data <= 5'd29;
94: data <= 5'd30;
95: data <= 5'd31;
96: data <= 5'd0;
97: data <= 5'd1;
98: data <= 5'd2;
99: data <= 5'd3;
100: data <= 5'd4;
101: data <= 5'd5;
102: data <= 5'd6;
103: data <= 5'd7;
104: data <= 5'd8;
105: data <= 5'd9;
106: data <= 5'd10;
107: data <= 5'd11;
108: data <= 5'd12;
109: data <= 5'd13;
110: data <= 5'd14;
111: data <= 5'd15;
112: data <= 5'd16;
113: data <= 5'd17;
114: data <= 5'd18;
115: data <= 5'd19;
116: data <= 5'd20;
117: data <= 5'd21;
118: data <= 5'd22;
119: data <= 5'd23;
120: data <= 5'd24;
121: data <= 5'd25;
122: data <= 5'd26;
123: data <= 5'd27;
124: data <= 5'd28;
125: data <= 5'd29;
126: data <= 5'd30;
127: data <= 5'd31;
    default : data <= 0;
    endcase
end
endmodule
