module mem_gen1 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 12;
input clk;
input [6:0] addr;
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= 12'd2285;
1: data <= 12'd872;
2: data <= 12'd1508;
3: data <= 12'd2333;
4: data <= 12'd3042;
5: data <= 12'd1779;
6: data <= 12'd282;
7: data <= 12'd1465;
8: data <= 12'd1602;
9: data <= 12'd602;
10: data <= 12'd247;
11: data <= 12'd870;
12: data <= 12'd1474;
13: data <= 12'd1755;
14: data <= 12'd3203;
15: data <= 12'd1187;
16: data <= 12'd205;
17: data <= 12'd156;
18: data <= 12'd2652;
19: data <= 12'd1807;
20: data <= 12'd758;
21: data <= 12'd2899;
22: data <= 12'd2677;
23: data <= 12'd2232;
24: data <= 12'd1325;
25: data <= 12'd2551;
26: data <= 12'd90;
27: data <= 12'd1530;
28: data <= 12'd2707;
29: data <= 12'd2742;
30: data <= 12'd8;
31: data <= 12'd136;
32: data <= 12'd2312;
33: data <= 12'd2685;
34: data <= 12'd2368;
35: data <= 12'd308;
36: data <= 12'd1907;
37: data <= 12'd2458;
38: data <= 12'd1838;
39: data <= 12'd1285;
40: data <= 12'd1871;
41: data <= 12'd1846;
42: data <= 12'd1421;
43: data <= 12'd854;
44: data <= 12'd1202;
45: data <= 12'd460;
46: data <= 12'd1162;
47: data <= 12'd3109;
48: data <= 12'd2918;
49: data <= 12'd3000;
50: data <= 12'd1065;
51: data <= 12'd1460;
52: data <= 12'd1517;
53: data <= 12'd2486;
54: data <= 12'd2314;
55: data <= 12'd2719;
56: data <= 12'd2946;
57: data <= 12'd147;
58: data <= 12'd2499;
59: data <= 12'd2535;
60: data <= 12'd3147;
61: data <= 12'd235;
62: data <= 12'd666;
63: data <= 12'd1335;
64: data <= 12'd2721;
65: data <= 12'd2980;
66: data <= 12'd725;
67: data <= 12'd2338;
68: data <= 12'd3127;
69: data <= 12'd3224;
70: data <= 12'd1544;
71: data <= 12'd2945;
72: data <= 12'd130;
73: data <= 12'd2210;
74: data <= 12'd951;
75: data <= 12'd2851;
76: data <= 12'd1861;
77: data <= 12'd1676;
78: data <= 12'd1860;
79: data <= 12'd1659;
80: data <= 12'd1571;
81: data <= 12'd75;
82: data <= 12'd1275;
83: data <= 12'd1701;
84: data <= 12'd2285;
85: data <= 12'd2226;
86: data <= 12'd1223;
87: data <= 12'd817;
88: data <= 12'd573;
89: data <= 12'd3083;
90: data <= 12'd2476;
91: data <= 12'd2144;
92: data <= 12'd3158;
93: data <= 12'd422;
94: data <= 12'd516;
95: data <= 12'd2114;
96: data <= 12'd2648;
97: data <= 12'd1739;
98: data <= 12'd2931;
99: data <= 12'd3221;
100: data <= 12'd1493;
101: data <= 12'd2078;
102: data <= 12'd2036;
103: data <= 12'd1322;
104: data <= 12'd2500;
105: data <= 12'd2552;
106: data <= 12'd107;
107: data <= 12'd1819;
108: data <= 12'd962;
109: data <= 12'd3038;
110: data <= 12'd1711;
111: data <= 12'd2455;
112: data <= 12'd1787;
113: data <= 12'd418;
114: data <= 12'd448;
115: data <= 12'd958;
116: data <= 12'd2970;
117: data <= 12'd555;
118: data <= 12'd2777;
119: data <= 12'd603;
120: data <= 12'd264;
121: data <= 12'd1159;
122: data <= 12'd3058;
123: data <= 12'd2051;
124: data <= 12'd1577;
125: data <= 12'd177;
126: data <= 12'd3009;
127: data <= 12'd1218;
    default : data <= 0;
    endcase
end
endmodule
