module tb_k2red;
