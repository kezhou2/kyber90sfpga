module mem_gen4 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 18;
input clk;
input [6:0] addr;//127
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= {6'd2,6'd1,6'd0};
1: data <= {6'd2,6'd1,6'd0};
2: data <= {6'd2,6'd1,6'd0};
3: data <= {6'd2,6'd1,6'd0};
4: data <= {6'd2,6'd1,6'd0};
5: data <= {6'd2,6'd1,6'd0};
6: data <= {6'd2,6'd1,6'd0};
7: data <= {6'd2,6'd1,6'd0};
8: data <= {6'd2,6'd1,6'd0};
9: data <= {6'd2,6'd1,6'd0};
10: data <= {6'd2,6'd1,6'd0};
11: data <= {6'd2,6'd1,6'd0};
12: data <= {6'd2,6'd1,6'd0};
13: data <= {6'd2,6'd1,6'd0};
14: data <= {6'd2,6'd1,6'd0};
15: data <= {6'd2,6'd1,6'd0};
16: data <= {6'd2,6'd1,6'd0};
17: data <= {6'd2,6'd1,6'd0};
18: data <= {6'd2,6'd1,6'd0};
19: data <= {6'd2,6'd1,6'd0};
20: data <= {6'd2,6'd1,6'd0};
21: data <= {6'd2,6'd1,6'd0};
22: data <= {6'd2,6'd1,6'd0};
23: data <= {6'd2,6'd1,6'd0};
24: data <= {6'd2,6'd1,6'd0};
25: data <= {6'd2,6'd1,6'd0};
26: data <= {6'd2,6'd1,6'd0};
27: data <= {6'd2,6'd1,6'd0};
28: data <= {6'd2,6'd1,6'd0};
29: data <= {6'd2,6'd1,6'd0};
30: data <= {6'd2,6'd1,6'd0};
31: data <= {6'd2,6'd1,6'd0};
32: data <= {6'd8,6'd7,6'd3};
33: data <= {6'd8,6'd7,6'd3};
34: data <= {6'd8,6'd7,6'd3};
35: data <= {6'd8,6'd7,6'd3};
36: data <= {6'd8,6'd7,6'd3};
37: data <= {6'd8,6'd7,6'd3};
38: data <= {6'd8,6'd7,6'd3};
39: data <= {6'd8,6'd7,6'd3};
40: data <= {6'd10,6'd9,6'd4};
41: data <= {6'd10,6'd9,6'd4};
42: data <= {6'd10,6'd9,6'd4};
43: data <= {6'd10,6'd9,6'd4};
44: data <= {6'd10,6'd9,6'd4};
45: data <= {6'd10,6'd9,6'd4};
46: data <= {6'd10,6'd9,6'd4};
47: data <= {6'd10,6'd9,6'd4};
48: data <= {6'd12,6'd11,6'd5};
49: data <= {6'd12,6'd11,6'd5};
50: data <= {6'd12,6'd11,6'd5};
51: data <= {6'd12,6'd11,6'd5};
52: data <= {6'd12,6'd11,6'd5};
53: data <= {6'd12,6'd11,6'd5};
54: data <= {6'd12,6'd11,6'd5};
55: data <= {6'd12,6'd11,6'd5};
56: data <= {6'd14,6'd13,6'd6};
57: data <= {6'd14,6'd13,6'd6};
58: data <= {6'd14,6'd13,6'd6};
59: data <= {6'd14,6'd13,6'd6};
60: data <= {6'd14,6'd13,6'd6};
61: data <= {6'd14,6'd13,6'd6};
62: data <= {6'd14,6'd13,6'd6};
63: data <= {6'd14,6'd13,6'd6};
64: data <= {6'd32,6'd31,6'd15};
65: data <= {6'd32,6'd31,6'd15};
66: data <= {6'd34,6'd33,6'd16};
67: data <= {6'd34,6'd33,6'd16};
68: data <= {6'd36,6'd35,6'd17};
69: data <= {6'd36,6'd35,6'd17};
70: data <= {6'd38,6'd37,6'd18};
71: data <= {6'd38,6'd37,6'd18};
72: data <= {6'd40,6'd39,6'd19};
73: data <= {6'd40,6'd39,6'd19};
74: data <= {6'd42,6'd41,6'd20};
75: data <= {6'd42,6'd41,6'd20};
76: data <= {6'd44,6'd43,6'd21};
77: data <= {6'd44,6'd43,6'd21};
78: data <= {6'd46,6'd45,6'd22};
79: data <= {6'd46,6'd45,6'd22};
80: data <= {6'd48,6'd47,6'd23};
81: data <= {6'd48,6'd47,6'd23};
82: data <= {6'd50,6'd49,6'd24};
83: data <= {6'd50,6'd49,6'd24};
84: data <= {6'd52,6'd51,6'd25};
85: data <= {6'd52,6'd51,6'd25};
86: data <= {6'd54,6'd53,6'd26};
87: data <= {6'd54,6'd53,6'd26};
88: data <= {6'd56,6'd55,6'd27};
89: data <= {6'd56,6'd55,6'd27};
90: data <= {6'd58,6'd57,6'd28};
91: data <= {6'd58,6'd57,6'd28};
92: data <= {6'd60,6'd59,6'd29};
93: data <= {6'd60,6'd59,6'd29};
94: data <= {6'd62,6'd61,6'd30};
95: data <= {6'd62,6'd61,6'd30};
96: data <= {6'd0,6'd4,6'd0};
97: data <= {6'd1,6'd5,6'd0};
98: data <= {6'd2,6'd6,6'd0};
99: data <= {6'd3,6'd7,6'd0};
100: data <= {6'd8,6'd12,6'd0};
101: data <= {6'd9,6'd13,6'd0};
102: data <= {6'd10,6'd14,6'd0};
103: data <= {6'd11,6'd15,6'd0};
104: data <= {6'd16,6'd20,6'd0};
105: data <= {6'd17,6'd21,6'd0};
106: data <= {6'd18,6'd22,6'd0};
107: data <= {6'd19,6'd23,6'd0};
108: data <= {6'd24,6'd28,6'd0};
109: data <= {6'd25,6'd29,6'd0};
110: data <= {6'd26,6'd30,6'd0};
111: data <= {6'd27,6'd31,6'd0};
112: data <= {6'd32,6'd36,6'd0};
113: data <= {6'd33,6'd37,6'd0};
114: data <= {6'd34,6'd38,6'd0};
115: data <= {6'd35,6'd39,6'd0};
116: data <= {6'd40,6'd44,6'd0};
117: data <= {6'd41,6'd45,6'd0};
118: data <= {6'd42,6'd46,6'd0};
119: data <= {6'd43,6'd47,6'd0};
120: data <= {6'd48,6'd52,6'd0};
121: data <= {6'd49,6'd53,6'd0};
122: data <= {6'd50,6'd54,6'd0};
123: data <= {6'd51,6'd55,6'd0};
124: data <= {6'd56,6'd60,6'd0};
125: data <= {6'd57,6'd61,6'd0};
126: data <= {6'd58,6'd62,6'd0};
127: data <= {6'd59,6'd63,6'd0};

    default : data <= 0;
    endcase
end
endmodule
