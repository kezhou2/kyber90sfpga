module mem_gen4 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 7*4;
input clk;
input [6:0] addr;//127
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= {7'd96,7'd32,7'd64,7'd64};
1: data <= {7'd96,7'd32,7'd64,7'd64};
2: data <= {7'd96,7'd32,7'd64,7'd64};
3: data <= {7'd96,7'd32,7'd64,7'd64};
4: data <= {7'd96,7'd32,7'd64,7'd64};
5: data <= {7'd96,7'd32,7'd64,7'd64};
6: data <= {7'd96,7'd32,7'd64,7'd64};
7: data <= {7'd96,7'd32,7'd64,7'd64};
8: data <= {7'd96,7'd32,7'd64,7'd64};
9: data <= {7'd96,7'd32,7'd64,7'd64};
10: data <= {7'd96,7'd32,7'd64,7'd64};
11: data <= {7'd96,7'd32,7'd64,7'd64};
12: data <= {7'd96,7'd32,7'd64,7'd64};
13: data <= {7'd96,7'd32,7'd64,7'd64};
14: data <= {7'd96,7'd32,7'd64,7'd64};
15: data <= {7'd96,7'd32,7'd64,7'd64};
16: data <= {7'd96,7'd32,7'd64,7'd64};
17: data <= {7'd96,7'd32,7'd64,7'd64};
18: data <= {7'd96,7'd32,7'd64,7'd64};
19: data <= {7'd96,7'd32,7'd64,7'd64};
20: data <= {7'd96,7'd32,7'd64,7'd64};
21: data <= {7'd96,7'd32,7'd64,7'd64};
22: data <= {7'd96,7'd32,7'd64,7'd64};
23: data <= {7'd96,7'd32,7'd64,7'd64};
24: data <= {7'd96,7'd32,7'd64,7'd64};
25: data <= {7'd96,7'd32,7'd64,7'd64};
26: data <= {7'd96,7'd32,7'd64,7'd64};
27: data <= {7'd96,7'd32,7'd64,7'd64};
28: data <= {7'd96,7'd32,7'd64,7'd64};
29: data <= {7'd96,7'd32,7'd64,7'd64};
30: data <= {7'd96,7'd32,7'd64,7'd64};
31: data <= {7'd96,7'd32,7'd64,7'd64};
32: data <= {7'd72,7'd8,7'd16,7'd16};
33: data <= {7'd72,7'd8,7'd16,7'd16};
34: data <= {7'd72,7'd8,7'd16,7'd16};
35: data <= {7'd72,7'd8,7'd16,7'd16};
36: data <= {7'd72,7'd8,7'd16,7'd16};
37: data <= {7'd72,7'd8,7'd16,7'd16};
38: data <= {7'd72,7'd8,7'd16,7'd16};
39: data <= {7'd72,7'd8,7'd16,7'd16};
40: data <= {7'd104,7'd40,7'd80,7'd80};
41: data <= {7'd104,7'd40,7'd80,7'd80};
42: data <= {7'd104,7'd40,7'd80,7'd80};
43: data <= {7'd104,7'd40,7'd80,7'd80};
44: data <= {7'd104,7'd40,7'd80,7'd80};
45: data <= {7'd104,7'd40,7'd80,7'd80};
46: data <= {7'd104,7'd40,7'd80,7'd80};
47: data <= {7'd104,7'd40,7'd80,7'd80};
48: data <= {7'd88,7'd24,7'd48,7'd48};
49: data <= {7'd88,7'd24,7'd48,7'd48};
50: data <= {7'd88,7'd24,7'd48,7'd48};
51: data <= {7'd88,7'd24,7'd48,7'd48};
52: data <= {7'd88,7'd24,7'd48,7'd48};
53: data <= {7'd88,7'd24,7'd48,7'd48};
54: data <= {7'd88,7'd24,7'd48,7'd48};
55: data <= {7'd88,7'd24,7'd48,7'd48};
56: data <= {7'd120,7'd56,7'd112,7'd112};
57: data <= {7'd120,7'd56,7'd112,7'd112};
58: data <= {7'd120,7'd56,7'd112,7'd112};
59: data <= {7'd120,7'd56,7'd112,7'd112};
60: data <= {7'd120,7'd56,7'd112,7'd112};
61: data <= {7'd120,7'd56,7'd112,7'd112};
62: data <= {7'd120,7'd56,7'd112,7'd112};
63: data <= {7'd120,7'd56,7'd112,7'd112};
64: data <= {7'd66,7'd2,7'd4,7'd4};
65: data <= {7'd66,7'd2,7'd4,7'd4};
66: data <= {7'd98,7'd34,7'd68,7'd68};
67: data <= {7'd98,7'd34,7'd68,7'd68};
68: data <= {7'd82,7'd18,7'd36,7'd36};
69: data <= {7'd82,7'd18,7'd36,7'd36};
70: data <= {7'd114,7'd50,7'd100,7'd100};
71: data <= {7'd114,7'd50,7'd100,7'd100};
72: data <= {7'd74,7'd10,7'd20,7'd20};
73: data <= {7'd74,7'd10,7'd20,7'd20};
74: data <= {7'd106,7'd42,7'd84,7'd84};
75: data <= {7'd106,7'd42,7'd84,7'd84};
76: data <= {7'd90,7'd26,7'd52,7'd52};
77: data <= {7'd90,7'd26,7'd52,7'd52};
78: data <= {7'd122,7'd58,7'd116,7'd116};
79: data <= {7'd122,7'd58,7'd116,7'd116};
80: data <= {7'd70,7'd6,7'd12,7'd12};
81: data <= {7'd70,7'd6,7'd12,7'd12};
82: data <= {7'd102,7'd38,7'd76,7'd76};
83: data <= {7'd102,7'd38,7'd76,7'd76};
84: data <= {7'd86,7'd22,7'd44,7'd44};
85: data <= {7'd86,7'd22,7'd44,7'd44};
86: data <= {7'd118,7'd54,7'd108,7'd108};
87: data <= {7'd118,7'd54,7'd108,7'd108};
88: data <= {7'd78,7'd14,7'd28,7'd28};
89: data <= {7'd78,7'd14,7'd28,7'd28};
90: data <= {7'd110,7'd46,7'd92,7'd92};
91: data <= {7'd110,7'd46,7'd92,7'd92};
92: data <= {7'd94,7'd30,7'd60,7'd60};
93: data <= {7'd94,7'd30,7'd60,7'd60};
94: data <= {7'd126,7'd62,7'd124,7'd124};
95: data <= {7'd126,7'd62,7'd124,7'd124};
96: data <= {7'd1,7'd9,7'd0,7'd0};
97: data <= {7'd3,7'd11,7'd0,7'd0};
98: data <= {7'd5,7'd13,7'd0,7'd0};
99: data <= {7'd7,7'd15,7'd0,7'd0};
100: data <= {7'd17,7'd25,7'd0,7'd0};
101: data <= {7'd19,7'd27,7'd0,7'd0};
102: data <= {7'd21,7'd29,7'd0,7'd0};
103: data <= {7'd23,7'd31,7'd0,7'd0};
104: data <= {7'd33,7'd41,7'd0,7'd0};
105: data <= {7'd35,7'd43,7'd0,7'd0};
106: data <= {7'd37,7'd45,7'd0,7'd0};
107: data <= {7'd39,7'd47,7'd0,7'd0};
108: data <= {7'd49,7'd57,7'd0,7'd0};
109: data <= {7'd51,7'd59,7'd0,7'd0};
110: data <= {7'd53,7'd61,7'd0,7'd0};
111: data <= {7'd55,7'd63,7'd0,7'd0};
112: data <= {7'd65,7'd73,7'd0,7'd0};
113: data <= {7'd67,7'd75,7'd0,7'd0};
114: data <= {7'd69,7'd77,7'd0,7'd0};
115: data <= {7'd71,7'd79,7'd0,7'd0};
116: data <= {7'd81,7'd89,7'd0,7'd0};
117: data <= {7'd83,7'd91,7'd0,7'd0};
118: data <= {7'd85,7'd93,7'd0,7'd0};
119: data <= {7'd87,7'd95,7'd0,7'd0};
120: data <= {7'd97,7'd105,7'd0,7'd0};
121: data <= {7'd99,7'd107,7'd0,7'd0};
122: data <= {7'd101,7'd109,7'd0,7'd0};
123: data <= {7'd103,7'd111,7'd0,7'd0};
124: data <= {7'd113,7'd121,7'd0,7'd0};
125: data <= {7'd115,7'd123,7'd0,7'd0};
126: data <= {7'd117,7'd125,7'd0,7'd0};
127: data <= {7'd119,7'd127,7'd0,7'd0};
    default : data <= 0;
    endcase
end
endmodule
