module mem_gen1 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 12;
input clk;
input [6:0] addr;
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= 12'd2285;
1: data <= 12'd872;
2: data <= 12'd2167;
3: data <= 12'd2144;
4: data <= 12'd1602;
5: data <= 12'd843;
6: data <= 12'd2931;
7: data <= 12'd1187;
8: data <= 12'd182;
9: data <= 12'd2552;
10: data <= 12'd2677;
11: data <= 12'd991;
12: data <= 12'd1787;
13: data <= 12'd2742;
14: data <= 12'd2378;
15: data <= 12'd603;
16: data <= 12'd1907;
17: data <= 12'd3254;
18: data <= 12'd3009;
19: data <= 12'd854;
20: data <= 12'd2756;
21: data <= 12'd1550;
22: data <= 12'd1065;
23: data <= 12'd1215;
24: data <= 12'd1855;
25: data <= 12'd147;
26: data <= 12'd1293;
27: data <= 12'd1522;
28: data <= 12'd2721;
29: data <= 12'd291;
30: data <= 12'd3239;
31: data <= 12'd2945;
32: data <= 12'd359;
33: data <= 12'd644;
34: data <= 12'd1860;
35: data <= 12'd1278;
36: data <= 12'd1458;
37: data <= 12'd2226;
38: data <= 12'd1508;
39: data <= 12'd220;
40: data <= 12'd3158;
41: data <= 12'd602;
42: data <= 12'd1015;
43: data <= 12'd3221;
44: data <= 12'd205;
45: data <= 12'd3094;
46: data <= 12'd107;
47: data <= 12'd2232;
48: data <= 12'd202;
49: data <= 12'd418;
50: data <= 12'd8;
51: data <= 12'd478;
52: data <= 12'd264;
53: data <= 12'd2458;
54: data <= 12'd2054;
55: data <= 12'd1218;
56: data <= 12'd1202;
57: data <= 12'd246;
58: data <= 12'd3047;
59: data <= 12'd1460;
60: data <= 12'd681;
61: data <= 12'd1574;
62: data <= 12'd2499;
63: data <= 12'd2007;
64: data <= 12'd2571;
65: data <= 12'd2980;
66: data <= 12'd1618;
67: data <= 12'd1799;
68: data <= 12'd130;
69: data <= 12'd2774;
70: data <= 12'd961;
71: data <= 12'd1659;
72: data <= 12'd1752;
73: data <= 12'd1483;
74: data <= 12'd1223;
75: data <= 12'd2333;
76: data <= 12'd411;
77: data <= 12'd422;
78: data <= 12'd247;
79: data <= 12'd610;
80: data <= 12'd1493;
81: data <= 12'd156;
82: data <= 12'd2663;
83: data <= 12'd1819;
84: data <= 12'd1325;
85: data <= 12'd105;
86: data <= 12'd448;
87: data <= 12'd136;
88: data <= 12'd1468;
89: data <= 12'd1159;
90: data <= 12'd1838;
91: data <= 12'd1628;
92: data <= 12'd732;
93: data <= 12'd460;
94: data <= 12'd853;
95: data <= 12'd1864;
96: data <= 12'd1517;
97: data <= 12'd1590;
98: data <= 12'd126;
99: data <= 12'd2535;
100: data <= 12'd829;
101: data <= 12'd430;
102: data <= 12'd725;
103: data <= 12'd874;
104: data <= 12'd622;
105: data <= 12'd2210;
106: data <= 12'd552;
107: data <= 12'd3021;
108: data <= 12'd1571;
109: data <= 12'd3152;
110: data <= 12'd1908;
111: data <= 12'd817;
112: data <= 12'd3042;
113: data <= 12'd329;
114: data <= 12'd516;
115: data <= 12'd870;
116: data <= 12'd383;
117: data <= 12'd2078;
118: data <= 12'd2652;
119: data <= 12'd1994;
120: data <= 12'd962;
121: data <= 12'd2551;
122: data <= 12'd1785;
123: data <= 12'd958;
124: data <= 12'd2312;
125: data <= 12'd1653;
126: data <= 12'd3058;
127: data <= 12'd1285;
    default : data <= 0;
    endcase
end
endmodule
