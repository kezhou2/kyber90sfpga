module mem_gen5 (clk, addr, wr_ena, data);
parameter DATA_WIDTH = 12;
input clk;
input [6:0] addr;
input wr_ena;
output [DATA_WIDTH-1:0] data;
reg [DATA_WIDTH-1:0] data;
always@(posedge clk) begin
 case (addr)
0: data <= 12'd2285;
1: data <= 12'd2044;
2: data <= 12'd1491;
3: data <= 12'd871;
4: data <= 12'd1422;
5: data <= 12'd3021;
6: data <= 12'd961;
7: data <= 12'd644;
8: data <= 12'd1017;
9: data <= 12'd3193;
10: data <= 12'd3321;
11: data <= 12'd587;
12: data <= 12'd622;
13: data <= 12'd1799;
14: data <= 12'd3239;
15: data <= 12'd778;
16: data <= 12'd2004;
17: data <= 12'd1097;
18: data <= 12'd652;
19: data <= 12'd430;
20: data <= 12'd2571;
21: data <= 12'd1522;
22: data <= 12'd677;
23: data <= 12'd3173;
24: data <= 12'd3124;
25: data <= 12'd2142;
26: data <= 12'd126;
27: data <= 12'd1574;
28: data <= 12'd1855;
29: data <= 12'd2459;
30: data <= 12'd3082;
31: data <= 12'd2727;
32: data <= 12'd1727;
33: data <= 12'd1864;
34: data <= 12'd3047;
35: data <= 12'd1550;
36: data <= 12'd287;
37: data <= 12'd996;
38: data <= 12'd1821;
39: data <= 12'd2457;
40: data <= 12'd732;
41: data <= 12'd1218;
42: data <= 12'd3009;
43: data <= 12'd177;
44: data <= 12'd1577;
45: data <= 12'd2051;
46: data <= 12'd3058;
47: data <= 12'd1159;
48: data <= 12'd264;
49: data <= 12'd603;
50: data <= 12'd2777;
51: data <= 12'd555;
52: data <= 12'd2970;
53: data <= 12'd958;
54: data <= 12'd448;
55: data <= 12'd418;
56: data <= 12'd1787;
57: data <= 12'd2455;
58: data <= 12'd1711;
59: data <= 12'd3038;
60: data <= 12'd962;
61: data <= 12'd1819;
62: data <= 12'd107;
63: data <= 12'd2552;
64: data <= 12'd2500;
65: data <= 12'd1322;
66: data <= 12'd2036;
67: data <= 12'd2078;
68: data <= 12'd1493;
69: data <= 12'd3221;
70: data <= 12'd2931;
71: data <= 12'd1739;
72: data <= 12'd2648;
73: data <= 12'd2114;
74: data <= 12'd516;
75: data <= 12'd422;
76: data <= 12'd3158;
77: data <= 12'd2144;
78: data <= 12'd2476;
79: data <= 12'd3083;
80: data <= 12'd573;
81: data <= 12'd817;
82: data <= 12'd1223;
83: data <= 12'd2226;
84: data <= 12'd2285;
85: data <= 12'd1701;
86: data <= 12'd1275;
87: data <= 12'd75;
88: data <= 12'd1571;
89: data <= 12'd1659;
90: data <= 12'd1860;
91: data <= 12'd1676;
92: data <= 12'd1861;
93: data <= 12'd2851;
94: data <= 12'd951;
95: data <= 12'd2210;
96: data <= 12'd130;
97: data <= 12'd2945;
98: data <= 12'd1544;
99: data <= 12'd3224;
100: data <= 12'd3127;
101: data <= 12'd2338;
102: data <= 12'd725;
103: data <= 12'd2980;
104: data <= 12'd2721;
105: data <= 12'd1335;
106: data <= 12'd666;
107: data <= 12'd235;
108: data <= 12'd3147;
109: data <= 12'd2535;
110: data <= 12'd2499;
111: data <= 12'd147;
112: data <= 12'd2946;
113: data <= 12'd2719;
114: data <= 12'd2314;
115: data <= 12'd2486;
116: data <= 12'd1517;
117: data <= 12'd1460;
118: data <= 12'd1065;
119: data <= 12'd3000;
120: data <= 12'd2918;
121: data <= 12'd3109;
122: data <= 12'd1162;
123: data <= 12'd460;
124: data <= 12'd1202;
125: data <= 12'd854;
126: data <= 12'd1421;
127: data <= 12'd1846;
    default : data <= 0;
    endcase
end
endmodule
